/*module tb();
	reg clk;
	wire [15:0]check_ra;
	
	processor proc (.clk(clk),.check_ra(check_ra));
	
	initial
		begin
			clk=1'b0;
			forever #5 clk=~clk;
		end
endmodule */
