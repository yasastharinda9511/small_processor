module R1_check(a_bus , out_r1);
	input [15:0] a_bus;
	output [15:0] out_r1;

	assign out_r1= a_bus;
endmodule